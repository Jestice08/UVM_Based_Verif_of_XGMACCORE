package mac_pkg;

	import uvm_pkg::*;
	
	`include "mac_env.sv"
	//`include "mac_interface.sv"
	//`include "mac_tb.sv"
	`include "mac_test.sv"
	//`include "mac_top.sv"
	`include "rst_agent.sv"
	`include "rst_driver.sv"
	`include "rst_monitor.sv"
	`include "rst_seq_item.sv"
	`include "rst_sequence.sv"
	`include "rx_agent.sv"
	`include "rx_monitor.sv"
	`include "scoreboard.sv"
	`include "seq_of_commands.sv"
	`include "tx_agent.sv"
	`include "tx_driver.sv"
	`include "tx_monitor.sv"
	`include "tx_sequence.sv"
	`include "virtual_sequencer.sv"
	`include "wb_agent.sv"
	`include "wb_driver.sv"
	`include "wb_monitor.sv"
	`include "wb_seq_item.sv"
	`include "wb_sequence.sv"
	
	
endpackage:mac_pkg
