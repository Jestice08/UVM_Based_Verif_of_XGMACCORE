//*********************************************
//          UVM Based Verification of         *
//           10 Gb Ethernet MAC Core          *
//                                            *
// Team member: Xuezhi Teng (xt2276)          *
//              Yi Zheng    (yz24299)         *
//*********************************************


// This is define file. It is used for defining some constants.

`define CPUREG_CONFIG0      8'h00
`define CPUREG_INT_PENDING  8'h08
`define CPUREG_INT_STATUS   8'h0c
`define CPUREG_INT_MASK     8'h10